i am in test
